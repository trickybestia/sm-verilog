// Port 1 - always read.
// Port 2 - read/write.

// Port 2 modes
`define MEM_READ       2'b00
`define MEM_WRITE_BYTE 2'b01
`define MEM_WRITE_HALF 2'b10
`define MEM_WRITE_WORD 2'b11
