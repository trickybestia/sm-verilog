typedef bit [15:0] UInt16;
typedef bit [3:0] Digit;

parameter EmptyDigit = 10;
