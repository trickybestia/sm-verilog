typedef bit [3:0] digit_t;

localparam empty_digit = 10;
