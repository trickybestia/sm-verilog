module AND1(input A, output Y);
    assign Y = A;
endmodule
